magic
tech sky130A
timestamp 1607430527
<< nwell >>
rect -17 185 722 315
<< nmos >>
rect 35 50 50 90
rect 150 75 165 115
rect 205 75 220 115
rect 320 75 335 115
rect 375 75 390 115
rect 485 75 500 115
rect 540 75 555 115
rect 655 50 670 90
<< pmos >>
rect 35 230 50 270
rect 150 205 165 245
rect 205 220 220 270
rect 320 205 335 245
rect 375 220 390 270
rect 485 220 500 270
rect 540 205 555 245
rect 655 230 670 270
<< ndiff >>
rect 116 105 150 115
rect 1 80 35 90
rect 1 60 5 80
rect 25 60 35 80
rect 1 50 35 60
rect 50 80 84 90
rect 50 60 60 80
rect 80 60 84 80
rect 116 85 120 105
rect 140 85 150 105
rect 116 75 150 85
rect 165 105 205 115
rect 165 85 175 105
rect 195 85 205 105
rect 165 75 205 85
rect 220 105 254 115
rect 220 85 230 105
rect 250 85 254 105
rect 220 75 254 85
rect 286 105 320 115
rect 286 85 290 105
rect 310 85 320 105
rect 286 75 320 85
rect 335 105 375 115
rect 335 85 345 105
rect 365 85 375 105
rect 335 75 375 85
rect 390 105 424 115
rect 390 85 400 105
rect 420 85 424 105
rect 390 75 424 85
rect 451 105 485 115
rect 451 85 455 105
rect 475 85 485 105
rect 451 75 485 85
rect 500 105 540 115
rect 500 85 510 105
rect 530 85 540 105
rect 500 75 540 85
rect 555 105 589 115
rect 555 85 565 105
rect 585 85 589 105
rect 555 75 589 85
rect 621 80 655 90
rect 50 50 84 60
rect 621 60 625 80
rect 645 60 655 80
rect 621 50 655 60
rect 670 80 704 90
rect 670 60 680 80
rect 700 60 704 80
rect 670 50 704 60
<< pdiff >>
rect 1 260 35 270
rect 1 240 5 260
rect 25 240 35 260
rect 1 230 35 240
rect 50 260 84 270
rect 50 240 60 260
rect 80 240 84 260
rect 50 230 84 240
rect 180 252 205 270
rect 178 250 205 252
rect 173 246 205 250
rect 173 245 178 246
rect 116 235 150 245
rect 116 215 120 235
rect 140 215 150 235
rect 116 205 150 215
rect 165 229 178 245
rect 195 229 205 246
rect 165 220 205 229
rect 220 260 254 270
rect 220 240 230 260
rect 250 240 254 260
rect 220 220 254 240
rect 165 205 190 220
rect 350 252 375 270
rect 348 250 375 252
rect 343 246 375 250
rect 343 245 348 246
rect 286 235 320 245
rect 286 215 290 235
rect 310 215 320 235
rect 286 205 320 215
rect 335 229 348 245
rect 365 229 375 246
rect 335 220 375 229
rect 390 260 424 270
rect 390 240 400 260
rect 420 240 424 260
rect 390 220 424 240
rect 451 260 485 270
rect 451 240 455 260
rect 475 240 485 260
rect 451 220 485 240
rect 500 252 525 270
rect 500 250 527 252
rect 500 246 532 250
rect 500 229 510 246
rect 527 245 532 246
rect 527 229 540 245
rect 500 220 540 229
rect 335 205 360 220
rect 515 205 540 220
rect 555 235 589 245
rect 555 215 565 235
rect 585 215 589 235
rect 555 205 589 215
rect 621 260 655 270
rect 621 240 625 260
rect 645 240 655 260
rect 621 230 655 240
rect 670 260 704 270
rect 670 240 680 260
rect 700 240 704 260
rect 670 230 704 240
<< ndiffc >>
rect 5 60 25 80
rect 60 60 80 80
rect 120 85 140 105
rect 175 85 195 105
rect 230 85 250 105
rect 290 85 310 105
rect 345 85 365 105
rect 400 85 420 105
rect 455 85 475 105
rect 510 85 530 105
rect 565 85 585 105
rect 625 60 645 80
rect 680 60 700 80
<< pdiffc >>
rect 5 240 25 260
rect 60 240 80 260
rect 120 215 140 235
rect 178 229 195 246
rect 230 240 250 260
rect 290 215 310 235
rect 348 229 365 246
rect 400 240 420 260
rect 455 240 475 260
rect 510 229 527 246
rect 565 215 585 235
rect 625 240 645 260
rect 680 240 700 260
<< poly >>
rect 35 270 50 284
rect 92 280 390 295
rect 35 183 50 230
rect 92 183 108 280
rect 205 270 220 280
rect 150 245 165 259
rect 205 206 220 220
rect 10 175 50 183
rect 10 155 15 175
rect 34 155 50 175
rect 10 147 50 155
rect 71 175 108 183
rect 150 195 165 205
rect 150 185 184 195
rect 150 180 220 185
rect 71 155 76 175
rect 95 155 108 175
rect 169 170 220 180
rect 71 147 108 155
rect 35 90 50 147
rect 92 145 108 147
rect 92 130 165 145
rect 150 115 165 130
rect 205 115 220 170
rect 262 145 278 280
rect 375 270 390 280
rect 485 280 613 295
rect 485 270 500 280
rect 320 245 335 259
rect 540 245 555 259
rect 375 206 390 220
rect 485 206 500 220
rect 320 195 335 205
rect 540 195 555 205
rect 320 185 354 195
rect 521 185 555 195
rect 320 180 390 185
rect 339 170 390 180
rect 262 130 335 145
rect 320 115 335 130
rect 375 115 390 170
rect 485 180 555 185
rect 597 183 613 280
rect 655 270 670 284
rect 655 183 670 230
rect 485 170 536 180
rect 597 175 634 183
rect 485 115 500 170
rect 597 155 610 175
rect 629 155 634 175
rect 597 147 634 155
rect 655 175 697 183
rect 655 155 670 175
rect 689 155 697 175
rect 655 147 697 155
rect 597 145 613 147
rect 540 130 613 145
rect 540 115 555 130
rect 655 90 670 147
rect 150 61 165 75
rect 35 40 50 50
rect 205 40 220 75
rect 320 61 335 75
rect 375 40 390 75
rect 35 25 390 40
rect 485 40 500 75
rect 540 61 555 75
rect 655 40 670 50
rect 485 25 670 40
<< polycont >>
rect 15 155 34 175
rect 76 155 95 175
rect 610 155 629 175
rect 670 155 689 175
<< locali >>
rect 5 260 25 285
rect 5 230 25 240
rect 60 260 80 280
rect 10 175 40 183
rect 10 155 15 175
rect 35 155 40 175
rect 10 147 40 155
rect 60 175 80 240
rect 120 235 140 270
rect 60 155 76 175
rect 95 155 103 175
rect 5 80 25 90
rect 5 35 25 60
rect 60 80 80 155
rect 120 105 140 215
rect 120 75 140 85
rect 175 246 195 270
rect 175 229 178 246
rect 175 190 195 229
rect 175 105 195 170
rect 175 75 195 85
rect 230 260 250 270
rect 230 105 250 240
rect 230 75 250 85
rect 290 235 310 270
rect 290 105 310 215
rect 290 75 310 85
rect 345 246 365 270
rect 345 229 348 246
rect 345 150 365 229
rect 345 105 365 130
rect 345 75 365 85
rect 400 260 420 270
rect 400 105 420 240
rect 400 75 420 85
rect 455 260 475 270
rect 455 150 475 240
rect 455 105 475 130
rect 455 75 475 85
rect 510 246 530 270
rect 527 229 530 246
rect 510 105 530 229
rect 510 75 530 85
rect 565 235 585 270
rect 565 190 585 215
rect 625 260 645 280
rect 625 175 645 240
rect 680 260 700 285
rect 680 230 700 240
rect 565 105 585 170
rect 602 155 610 175
rect 629 155 645 175
rect 565 75 585 85
rect 625 80 645 155
rect 665 175 695 183
rect 665 155 670 175
rect 690 155 695 175
rect 665 147 695 155
rect 60 50 80 60
rect 625 50 645 60
rect 680 80 700 90
rect 680 35 700 60
<< viali >>
rect 5 285 25 305
rect 680 285 700 305
rect 15 155 34 175
rect 34 155 35 175
rect 175 170 195 190
rect 345 130 365 150
rect 455 130 475 150
rect 565 170 585 190
rect 670 155 689 175
rect 689 155 690 175
rect 5 15 25 35
rect 680 15 700 35
<< metal1 >>
rect 1 305 704 320
rect 1 285 5 305
rect 25 285 680 305
rect 700 285 704 305
rect 1 270 704 285
rect 170 190 200 195
rect 560 190 590 195
rect 8 175 42 183
rect 8 155 15 175
rect 35 155 42 175
rect 169 170 175 190
rect 195 170 565 190
rect 585 170 591 190
rect 663 175 697 183
rect 170 165 200 170
rect 560 165 590 170
rect 663 155 670 175
rect 690 155 697 175
rect 8 147 42 155
rect 340 150 370 155
rect 450 150 480 155
rect 339 130 345 150
rect 365 130 455 150
rect 475 130 481 150
rect 663 147 697 155
rect 340 125 370 130
rect 450 125 480 130
rect 1 35 705 50
rect 1 15 5 35
rect 25 15 680 35
rect 700 15 705 35
rect 1 0 705 15
<< end >>
