///////// CARRY CHAIN /////////

module clb #() ();

endmodule
