magic
tech sky130A
timestamp 1607344602
<< nwell >>
rect -15 190 775 315
rect -15 185 120 190
rect 262 185 775 190
<< nmos >>
rect 40 50 55 90
rect 155 50 170 90
rect 210 50 225 90
rect 345 50 360 90
rect 400 50 415 90
rect 540 50 555 90
rect 595 50 610 90
rect 705 50 720 90
<< pmos >>
rect 40 230 55 270
rect 155 230 170 270
rect 210 230 225 270
rect 345 230 360 270
rect 400 230 415 270
rect 540 230 555 270
rect 595 230 610 270
rect 705 230 720 270
<< ndiff >>
rect 5 80 40 90
rect 5 60 10 80
rect 30 60 40 80
rect 5 50 40 60
rect 55 80 90 90
rect 55 60 65 80
rect 85 60 90 80
rect 55 50 90 60
rect 120 80 155 90
rect 120 60 125 80
rect 145 60 155 80
rect 120 50 155 60
rect 170 80 210 90
rect 170 60 180 80
rect 200 60 210 80
rect 170 50 210 60
rect 225 80 260 90
rect 225 60 235 80
rect 255 60 260 80
rect 225 50 260 60
rect 310 80 345 90
rect 310 60 315 80
rect 335 60 345 80
rect 310 50 345 60
rect 360 80 400 90
rect 360 60 370 80
rect 390 60 400 80
rect 360 50 400 60
rect 415 80 450 90
rect 415 60 425 80
rect 445 60 450 80
rect 415 50 450 60
rect 505 80 540 90
rect 505 60 510 80
rect 530 60 540 80
rect 505 50 540 60
rect 555 80 595 90
rect 555 60 565 80
rect 585 60 595 80
rect 555 50 595 60
rect 610 80 644 90
rect 610 60 620 80
rect 640 60 644 80
rect 610 50 644 60
rect 671 80 705 90
rect 671 60 675 80
rect 695 60 705 80
rect 671 50 705 60
rect 720 80 755 90
rect 720 60 730 80
rect 750 60 755 80
rect 720 50 755 60
<< pdiff >>
rect 5 260 40 270
rect 5 240 10 260
rect 30 240 40 260
rect 5 230 40 240
rect 55 260 89 270
rect 55 240 65 260
rect 85 240 89 260
rect 55 230 89 240
rect 121 260 155 270
rect 121 240 125 260
rect 145 240 155 260
rect 121 230 155 240
rect 170 260 210 270
rect 170 240 180 260
rect 200 240 210 260
rect 170 230 210 240
rect 225 260 260 270
rect 225 240 235 260
rect 255 240 260 260
rect 225 230 260 240
rect 311 260 345 270
rect 311 240 315 260
rect 335 240 345 260
rect 311 230 345 240
rect 360 260 400 270
rect 360 240 370 260
rect 390 240 400 260
rect 360 230 400 240
rect 415 260 449 270
rect 415 240 425 260
rect 445 240 449 260
rect 415 230 449 240
rect 506 260 540 270
rect 506 240 510 260
rect 530 240 540 260
rect 506 230 540 240
rect 555 260 595 270
rect 555 240 565 260
rect 585 240 595 260
rect 555 230 595 240
rect 610 260 644 270
rect 610 240 620 260
rect 640 240 644 260
rect 610 230 644 240
rect 671 260 705 270
rect 671 240 675 260
rect 695 240 705 260
rect 671 230 705 240
rect 720 260 755 270
rect 720 240 730 260
rect 750 240 755 260
rect 720 230 755 240
<< ndiffc >>
rect 10 60 30 80
rect 65 60 85 80
rect 125 60 145 80
rect 180 60 200 80
rect 235 60 255 80
rect 315 60 335 80
rect 370 60 390 80
rect 425 60 445 80
rect 510 60 530 80
rect 565 60 585 80
rect 620 60 640 80
rect 675 60 695 80
rect 730 60 750 80
<< pdiffc >>
rect 10 240 30 260
rect 65 240 85 260
rect 125 240 145 260
rect 180 240 200 260
rect 235 240 255 260
rect 315 240 335 260
rect 370 240 390 260
rect 425 240 445 260
rect 510 240 530 260
rect 565 240 585 260
rect 620 240 640 260
rect 675 240 695 260
rect 730 240 750 260
<< poly >>
rect 80 312 415 320
rect 80 295 86 312
rect 103 305 415 312
rect 103 295 108 305
rect 80 285 108 295
rect 40 270 55 285
rect 155 270 170 283
rect 210 270 225 305
rect 345 270 360 283
rect 400 270 415 305
rect 540 312 684 320
rect 540 305 657 312
rect 540 270 555 305
rect 648 295 657 305
rect 674 295 684 312
rect 648 290 679 295
rect 595 270 610 284
rect 705 270 720 284
rect 40 195 55 230
rect 155 210 170 230
rect 120 205 170 210
rect 120 195 130 205
rect 40 185 130 195
rect 150 185 170 205
rect 40 180 170 185
rect 40 90 55 180
rect 155 90 170 180
rect 210 90 225 230
rect 345 210 360 230
rect 310 205 360 210
rect 310 185 320 205
rect 340 185 360 205
rect 310 180 360 185
rect 345 90 360 180
rect 400 90 415 230
rect 540 206 555 230
rect 475 191 555 206
rect 40 35 55 50
rect 155 35 170 50
rect 210 35 225 50
rect 345 35 360 50
rect 400 35 415 50
rect 475 15 490 191
rect 595 170 610 230
rect 705 170 720 230
rect 540 155 720 170
rect 540 90 555 155
rect 595 90 610 105
rect 705 90 720 155
rect 540 36 555 50
rect 595 15 610 50
rect 705 35 720 50
rect 475 0 610 15
<< polycont >>
rect 86 295 103 312
rect 657 295 674 312
rect 130 185 150 205
rect 320 185 340 205
<< locali >>
rect 65 312 108 320
rect 10 260 30 285
rect 10 230 30 240
rect 65 295 86 312
rect 103 295 108 312
rect 648 312 695 320
rect 65 285 108 295
rect 125 290 295 310
rect 65 260 85 285
rect 10 80 30 90
rect 10 35 30 60
rect 65 80 85 240
rect 125 260 145 290
rect 125 230 145 240
rect 180 260 200 270
rect 125 205 155 210
rect 122 185 130 205
rect 150 185 160 205
rect 125 180 155 185
rect 180 165 200 240
rect 65 50 85 60
rect 125 80 145 110
rect 125 50 145 60
rect 180 80 200 145
rect 235 260 255 270
rect 235 130 255 240
rect 254 111 255 130
rect 235 110 255 111
rect 275 90 295 290
rect 315 290 485 310
rect 648 295 657 312
rect 674 295 695 312
rect 648 290 695 295
rect 315 260 335 290
rect 315 230 335 240
rect 370 260 390 270
rect 315 205 345 210
rect 370 205 390 240
rect 312 185 320 205
rect 340 185 350 205
rect 315 180 345 185
rect 180 50 200 60
rect 235 80 295 90
rect 255 70 295 80
rect 315 80 335 110
rect 235 50 255 60
rect 315 50 335 60
rect 370 80 390 185
rect 425 260 445 270
rect 425 130 445 240
rect 444 111 445 130
rect 425 110 445 111
rect 465 90 485 290
rect 370 50 390 60
rect 425 80 485 90
rect 445 70 485 80
rect 510 260 530 270
rect 510 205 530 240
rect 510 80 530 185
rect 425 50 445 60
rect 510 50 530 60
rect 565 260 585 270
rect 565 80 585 240
rect 565 50 585 60
rect 620 260 640 270
rect 620 170 640 240
rect 620 80 640 150
rect 620 50 640 60
rect 675 260 695 290
rect 675 80 695 240
rect 730 260 750 285
rect 730 230 750 240
rect 675 50 695 60
rect 730 80 750 90
rect 730 35 750 60
<< viali >>
rect 10 285 30 305
rect 130 185 150 205
rect 180 145 200 165
rect 125 110 145 130
rect 235 111 254 130
rect 320 185 340 205
rect 370 185 390 205
rect 315 110 335 130
rect 425 111 444 130
rect 510 185 530 205
rect 620 150 640 170
rect 730 285 750 305
rect 10 15 30 35
rect 730 15 750 35
<< metal1 >>
rect 5 305 755 320
rect 5 285 10 305
rect 30 285 730 305
rect 750 285 755 305
rect 5 270 755 285
rect 125 205 155 210
rect 315 205 345 210
rect 365 205 395 210
rect 505 205 535 210
rect 124 185 130 205
rect 150 185 320 205
rect 340 185 350 205
rect 364 185 370 205
rect 390 185 510 205
rect 530 185 536 205
rect 125 180 155 185
rect 315 180 345 185
rect 365 180 395 185
rect 505 180 535 185
rect 615 170 645 175
rect 175 165 205 170
rect 610 165 620 170
rect 174 145 180 165
rect 200 150 620 165
rect 640 150 646 170
rect 200 145 210 150
rect 615 145 645 150
rect 175 140 205 145
rect 120 130 150 135
rect 230 130 260 135
rect 310 130 340 135
rect 420 130 450 135
rect 119 110 125 130
rect 145 125 155 130
rect 225 125 235 130
rect 145 111 235 125
rect 254 111 261 130
rect 145 110 261 111
rect 309 110 315 130
rect 335 111 425 130
rect 444 111 451 130
rect 335 110 451 111
rect 120 105 150 110
rect 230 105 260 110
rect 310 105 340 110
rect 420 105 450 110
rect 5 35 755 50
rect 5 15 10 35
rect 30 15 730 35
rect 750 15 755 35
rect 5 0 755 15
<< labels >>
rlabel poly 40 145 55 180 1 S1
rlabel pdiffc 125 240 145 260 1 C
rlabel pdiffc 235 240 255 260 1 A
rlabel pdiffc 315 240 335 260 1 C
rlabel pdiffc 425 240 445 260 1 A
rlabel pdiffc 620 240 640 260 1 A
rlabel pdiffc 510 240 530 260 1 C
rlabel viali 12 18 27 32 1 VGND
rlabel viali 12 288 28 303 1 VPWR
rlabel poly 705 105 720 125 1 S2
rlabel locali 565 115 585 130 1 OUT
rlabel ndiffc 315 60 335 80 1 D
rlabel ndiffc 425 60 445 80 1 C
rlabel ndiffc 235 60 255 80 1 A
rlabel ndiffc 125 60 145 80 1 B
<< end >>
