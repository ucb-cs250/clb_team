magic
tech sky130A
timestamp 1607304229
<< nwell >>
rect -15 200 260 315
<< nmos >>
rect 40 50 55 90
rect 155 50 170 90
<< pmos >>
rect 40 230 55 270
rect 155 230 170 270
<< ndiff >>
rect 5 80 40 90
rect 5 60 10 80
rect 30 60 40 80
rect 5 50 40 60
rect 55 80 90 90
rect 55 60 65 80
rect 85 60 90 80
rect 55 50 90 60
rect 120 80 155 90
rect 120 60 125 80
rect 145 60 155 80
rect 120 50 155 60
rect 170 80 240 90
rect 170 60 180 80
rect 200 60 240 80
rect 170 50 240 60
<< pdiff >>
rect 5 260 40 270
rect 5 240 10 260
rect 30 240 40 260
rect 5 230 40 240
rect 55 260 90 270
rect 55 240 65 260
rect 85 240 90 260
rect 55 230 90 240
rect 120 260 155 270
rect 120 240 125 260
rect 145 240 155 260
rect 120 230 155 240
rect 170 260 240 270
rect 170 240 180 260
rect 200 240 240 260
rect 170 230 240 240
<< ndiffc >>
rect 10 60 30 80
rect 65 60 85 80
rect 125 60 145 80
rect 180 60 200 80
<< pdiffc >>
rect 10 240 30 260
rect 65 240 85 260
rect 125 240 145 260
rect 180 240 200 260
<< poly >>
rect 40 270 55 290
rect 155 270 170 290
rect 40 120 55 230
rect 95 200 125 205
rect 155 200 170 230
rect 90 180 100 200
rect 120 180 170 200
rect 95 175 125 180
rect 40 105 170 120
rect 40 90 55 105
rect 155 90 170 105
rect 40 30 55 50
rect 155 30 170 50
<< polycont >>
rect 100 180 120 200
<< locali >>
rect 10 260 30 285
rect 10 230 30 240
rect 65 260 85 270
rect 65 205 85 240
rect 125 260 145 270
rect 125 230 145 240
rect 180 260 200 270
rect 65 200 125 205
rect 65 180 100 200
rect 120 180 130 200
rect 65 175 125 180
rect 10 80 30 90
rect 10 35 30 60
rect 65 80 85 175
rect 65 50 85 60
rect 125 80 145 90
rect 125 50 145 60
rect 180 80 200 240
rect 180 50 200 60
<< viali >>
rect 10 285 30 305
rect 10 15 30 35
<< metal1 >>
rect 5 305 220 320
rect 5 285 10 305
rect 30 285 220 305
rect 5 270 220 285
rect 5 35 180 50
rect 5 15 10 35
rect 30 15 180 35
rect 5 0 180 15
<< end >>
