VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mux4i
  CLASS BLOCK ;
  FOREIGN mux4i ;
  ORIGIN 0.170 0.000 ;
  SIZE 7.940 BY 3.200 ;
  OBS
      LAYER nwell ;
        RECT -0.170 1.850 7.770 3.150 ;
      LAYER li1 ;
        RECT 0.050 2.300 0.250 3.050 ;
        RECT 0.100 1.470 0.400 1.830 ;
        RECT 0.600 1.750 0.800 2.800 ;
        RECT 0.600 1.550 1.030 1.750 ;
        RECT 0.050 0.150 0.250 0.900 ;
        RECT 0.600 0.500 0.800 1.550 ;
        RECT 1.200 0.750 1.400 2.700 ;
        RECT 1.750 0.750 1.950 2.700 ;
        RECT 2.300 0.750 2.500 2.700 ;
        RECT 2.900 0.750 3.100 2.700 ;
        RECT 3.450 0.750 3.650 2.700 ;
        RECT 4.000 0.750 4.200 2.700 ;
        RECT 4.550 0.750 4.750 2.700 ;
        RECT 5.100 0.750 5.300 2.700 ;
        RECT 5.650 0.750 5.850 2.700 ;
        RECT 6.250 1.750 6.450 2.800 ;
        RECT 6.800 2.320 7.000 3.050 ;
        RECT 6.620 1.790 6.920 2.150 ;
        RECT 6.020 1.550 6.450 1.750 ;
        RECT 6.250 0.500 6.450 1.550 ;
        RECT 6.880 1.220 7.180 1.580 ;
        RECT 7.350 1.500 7.550 2.800 ;
        RECT 7.350 1.300 7.600 1.500 ;
        RECT 6.800 0.150 7.000 0.900 ;
        RECT 7.350 0.400 7.550 1.300 ;
      LAYER mcon ;
        RECT 0.050 2.850 0.250 3.050 ;
        RECT 6.800 2.850 7.000 3.050 ;
        RECT 0.150 1.550 0.350 1.750 ;
        RECT 1.200 2.150 1.400 2.350 ;
        RECT 1.750 1.700 1.950 1.900 ;
        RECT 2.300 0.850 2.500 1.050 ;
        RECT 2.900 2.150 3.100 2.350 ;
        RECT 3.450 1.300 3.650 1.500 ;
        RECT 4.000 0.850 4.200 1.050 ;
        RECT 4.550 1.300 4.750 1.500 ;
        RECT 5.100 1.300 5.300 1.500 ;
        RECT 5.650 1.700 5.850 1.900 ;
        RECT 6.670 1.870 6.870 2.070 ;
        RECT 6.930 1.300 7.130 1.500 ;
        RECT 7.400 1.300 7.600 1.500 ;
      LAYER met1 ;
        RECT 0.010 2.700 7.590 3.200 ;
        RECT 1.150 2.360 1.450 2.400 ;
        RECT 1.140 2.150 1.460 2.360 ;
        RECT 2.850 2.350 3.160 2.400 ;
        RECT 2.840 2.150 3.160 2.350 ;
        RECT 1.150 2.100 1.450 2.150 ;
        RECT 2.850 2.100 3.160 2.150 ;
        RECT 1.700 1.900 2.000 1.950 ;
        RECT 5.600 1.900 5.900 1.950 ;
        RECT 0.080 1.470 0.420 1.830 ;
        RECT 1.690 1.700 5.910 1.900 ;
        RECT 6.600 1.790 6.940 2.150 ;
        RECT 1.700 1.650 2.000 1.700 ;
        RECT 5.600 1.650 5.900 1.700 ;
        RECT 3.400 1.500 3.700 1.550 ;
        RECT 4.500 1.500 4.800 1.550 ;
        RECT 5.050 1.500 5.350 1.550 ;
        RECT 6.860 1.500 7.200 1.580 ;
        RECT 7.350 1.500 7.650 1.550 ;
        RECT 3.390 1.300 4.810 1.500 ;
        RECT 5.040 1.300 7.200 1.500 ;
        RECT 7.340 1.300 7.660 1.500 ;
        RECT 3.400 1.250 3.700 1.300 ;
        RECT 4.500 1.250 4.800 1.300 ;
        RECT 5.050 1.250 5.350 1.300 ;
        RECT 6.860 1.220 7.200 1.300 ;
        RECT 7.350 1.250 7.650 1.300 ;
        RECT 2.250 1.050 2.550 1.100 ;
        RECT 3.950 1.050 4.250 1.100 ;
        RECT 2.240 0.850 2.560 1.050 ;
        RECT 3.940 0.850 4.260 1.050 ;
        RECT 2.250 0.800 2.550 0.850 ;
        RECT 3.950 0.800 4.250 0.850 ;
        RECT 0.010 0.000 7.590 0.500 ;
  END
END mux4i
END LIBRARY

