magic
tech sky130A
timestamp 1607334395
<< nwell >>
rect -15 185 320 315
<< nmos >>
rect 40 50 55 90
rect 155 50 170 90
rect 210 50 225 90
<< pmos >>
rect 40 230 55 270
rect 155 205 170 270
rect 210 205 225 270
<< ndiff >>
rect 5 80 40 90
rect 5 60 10 80
rect 30 60 40 80
rect 5 50 40 60
rect 55 80 90 90
rect 55 60 65 80
rect 85 60 90 80
rect 55 50 90 60
rect 120 80 155 90
rect 120 60 125 80
rect 145 60 155 80
rect 120 50 155 60
rect 170 80 210 90
rect 170 60 180 80
rect 200 60 210 80
rect 170 50 210 60
rect 225 80 300 90
rect 225 60 235 80
rect 255 60 300 80
rect 225 50 300 60
<< pdiff >>
rect 5 260 40 270
rect 5 240 10 260
rect 30 240 40 260
rect 5 230 40 240
rect 55 260 89 270
rect 55 240 65 260
rect 85 240 89 260
rect 55 230 89 240
rect 121 260 155 270
rect 121 240 125 260
rect 145 240 155 260
rect 121 205 155 240
rect 170 230 210 270
rect 170 210 180 230
rect 200 210 210 230
rect 170 205 210 210
rect 225 260 300 270
rect 225 240 235 260
rect 255 240 300 260
rect 225 205 300 240
<< ndiffc >>
rect 10 60 30 80
rect 65 60 85 80
rect 125 60 145 80
rect 180 60 200 80
rect 235 60 255 80
<< pdiffc >>
rect 10 240 30 260
rect 65 240 85 260
rect 125 240 145 260
rect 180 210 200 230
rect 235 240 255 260
<< poly >>
rect 80 312 225 320
rect 80 295 86 312
rect 103 305 225 312
rect 103 295 108 305
rect 80 285 108 295
rect 40 270 55 285
rect 155 270 170 283
rect 210 270 225 305
rect 40 195 55 230
rect 155 195 170 205
rect 40 180 170 195
rect 40 90 55 180
rect 155 90 170 180
rect 210 90 225 205
rect 40 35 55 50
rect 155 35 170 50
rect 210 35 225 50
<< polycont >>
rect 86 295 103 312
<< locali >>
rect 65 312 108 320
rect 10 260 30 285
rect 10 230 30 240
rect 65 295 86 312
rect 103 295 108 312
rect 65 285 108 295
rect 125 290 295 310
rect 65 260 85 285
rect 10 80 30 90
rect 10 35 30 60
rect 65 80 85 240
rect 125 260 145 290
rect 235 260 255 270
rect 125 225 145 240
rect 180 230 200 240
rect 65 50 85 60
rect 125 80 145 110
rect 125 50 145 60
rect 180 80 200 210
rect 235 130 255 240
rect 254 111 255 130
rect 235 110 255 111
rect 275 90 295 290
rect 180 50 200 60
rect 235 80 295 90
rect 255 70 295 80
rect 235 50 255 60
<< viali >>
rect 10 285 30 305
rect 125 110 145 130
rect 235 111 254 130
rect 10 15 30 35
<< metal1 >>
rect 5 305 300 320
rect 5 285 10 305
rect 30 285 300 305
rect 5 270 300 285
rect 120 130 150 135
rect 230 130 260 135
rect 119 110 125 130
rect 145 111 235 130
rect 254 111 261 130
rect 145 110 261 111
rect 120 105 150 110
rect 230 105 260 110
rect 5 48 275 50
rect 5 35 300 48
rect 5 15 10 35
rect 30 15 300 35
rect 5 0 300 15
<< labels >>
rlabel poly 40 145 55 180 1 S1
rlabel locali 185 135 195 155 1 out_AC
rlabel pdiffc 125 240 145 260 1 C
rlabel pdiffc 235 240 255 260 1 A
<< end >>
